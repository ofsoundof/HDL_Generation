module div_16bit (
    input wire [15:0] A,
    input wire [7:0] B,
    output reg [15:0] result,
    output reg [15:0] odd
);

reg [15:0] a_reg;
reg [7:0] b_reg;

always @(A or B) begin
    a_reg <= A;
    b_reg <= B;
end

always @(*) begin
    if (b_reg == 0) begin
        result = 0;
        odd = a_reg;
    end else begin
        reg [15:0] temp_result = 0;
        reg [15:0] temp_odd = a_reg;
        for (int i = 7; i >= 0; i = i - 1) begin
            if ((temp_odd << i) >= b_reg) begin
                temp_result[i] <= 1;
                temp_odd = temp_odd - (b_reg << i);
            end else begin
                temp_result[i] <= 0;
            end
        end
        result = temp_result;
        odd = temp_odd;
    end
end

endmodule